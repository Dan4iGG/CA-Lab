<<<<<<< HEAD
module ex1 (sw0, sw1, led0);
	input sw0, sw1;
	output led0;
	and (led0, sw0, sw1);
endmodule
=======
module ex1 (sw0, sw1, led0);
	input sw0, sw1;
	output led0;
	and (led0, sw0, sw1);
endmodule
>>>>>>> 4dcf63ba51e4d922f9c1cc83d9d3efef3a8f546f
